`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:49:25 09/05/2018 
// Design Name: 
// Module Name:    seven_seg_decoder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module seven_seg_decoder(bcd, blank, seg);
	input [3:0] bcd;
	input blank;
	output [7:1] seg;
	
	


endmodule
